magic
tech scmos
timestamp 1619529522
<< metal1 >>
rect 10 154 17 187
rect -108 46 -101 148
rect 35 139 42 187
rect 501 154 508 187
rect -96 85 -89 133
rect 165 -66 172 69
rect 181 24 188 133
rect 202 61 209 148
rect 354 -66 361 64
rect 383 46 390 148
rect 526 139 533 187
rect 992 154 999 187
rect 395 85 402 133
rect 656 -66 663 69
rect 672 24 679 133
rect 693 61 700 148
rect 845 -66 852 64
rect 874 51 881 148
rect 1017 139 1024 187
rect 1483 154 1490 187
rect 886 90 893 133
rect 1147 -66 1154 69
rect 1163 29 1170 133
rect 1184 67 1191 148
rect 1336 -66 1343 64
rect 1365 51 1372 148
rect 1509 139 1516 187
rect 1377 90 1384 133
rect 1638 -66 1645 69
rect 1654 29 1661 133
rect 1675 67 1682 148
rect 1827 -66 1834 64
<< m2contact >>
rect -108 148 -101 154
rect 10 148 17 154
rect 202 148 209 154
rect -96 133 -89 139
rect 35 133 42 139
rect 181 133 188 139
rect 96 122 103 128
rect 96 0 103 5
rect 383 148 390 154
rect 501 148 508 154
rect 220 122 227 128
rect 300 122 307 128
rect 223 0 230 5
rect 306 0 313 5
rect 693 148 700 154
rect 395 133 402 139
rect 526 133 533 139
rect 672 133 679 139
rect 419 122 426 128
rect 587 122 594 128
rect 435 0 442 5
rect 587 0 594 5
rect 874 148 881 154
rect 992 148 999 154
rect 711 122 718 128
rect 791 122 798 128
rect 714 0 721 5
rect 797 0 804 5
rect 1184 148 1191 154
rect 886 133 893 139
rect 1017 133 1024 139
rect 1163 133 1170 139
rect 910 122 917 128
rect 1078 122 1085 128
rect 926 0 933 5
rect 1078 0 1085 5
rect 1365 148 1372 154
rect 1483 148 1490 154
rect 1202 122 1209 128
rect 1282 122 1289 128
rect 1205 0 1212 5
rect 1288 0 1295 5
rect 1675 148 1682 154
rect 1377 133 1384 139
rect 1509 133 1516 139
rect 1654 133 1661 139
rect 1401 122 1408 128
rect 1569 122 1576 128
rect 1417 0 1424 5
rect 1569 0 1576 5
rect 1693 122 1700 128
rect 1696 0 1703 5
<< metal2 >>
rect -101 148 10 154
rect 17 148 202 154
rect 390 148 501 154
rect 508 148 693 154
rect 881 148 992 154
rect 999 148 1184 154
rect 1372 148 1483 154
rect 1490 148 1675 154
rect -89 133 35 139
rect 42 133 181 139
rect 402 133 526 139
rect 533 133 672 139
rect 893 133 1017 139
rect 1024 133 1163 139
rect 1384 133 1509 139
rect 1516 133 1654 139
rect 103 122 220 128
rect 307 122 419 128
rect 594 122 711 128
rect 798 122 910 128
rect 1085 122 1202 128
rect 1289 122 1401 128
rect 1576 122 1693 128
rect 103 0 223 5
rect 313 0 435 5
rect 594 0 714 5
rect 804 0 926 5
rect 1085 0 1205 5
rect 1295 0 1417 5
rect 1576 0 1696 5
use xorgate  xorgate_0
timestamp 1618846832
transform 1 0 34 0 1 53
box -142 -53 138 75
use andgate  andgate_0
timestamp 1618893190
transform 1 0 296 0 1 36
box -115 -36 65 92
use xorgate  xorgate_1
timestamp 1618846832
transform 1 0 525 0 1 53
box -142 -53 138 75
use andgate  andgate_1
timestamp 1618893190
transform 1 0 787 0 1 36
box -115 -36 65 92
use xorgate  xorgate_2
timestamp 1618846832
transform 1 0 1016 0 1 53
box -142 -53 138 75
use andgate  andgate_2
timestamp 1618893190
transform 1 0 1278 0 1 36
box -115 -36 65 92
use xorgate  xorgate_3
timestamp 1618846832
transform 1 0 1507 0 1 53
box -142 -53 138 75
use andgate  andgate_3
timestamp 1618893190
transform 1 0 1769 0 1 36
box -115 -36 65 92
<< end >>
