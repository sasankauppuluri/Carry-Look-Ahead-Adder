magic
tech scmos
timestamp 1619544759
<< metal1 >>
rect 196 1935 379 1942
rect 198 1746 361 1753
rect 0 1617 48 1624
rect 0 1591 33 1598
rect 253 1444 343 1451
rect 252 1255 325 1262
rect 316 1158 325 1255
rect 316 1153 320 1158
rect 0 1125 48 1132
rect 0 1100 33 1107
rect 253 953 307 960
rect 248 764 280 771
rect 0 634 48 641
rect 0 609 33 616
rect 235 462 271 469
rect 206 273 240 280
rect 0 143 48 150
rect 0 118 33 125
rect 244 62 253 273
rect 262 133 271 462
rect 280 223 289 764
rect 298 322 307 953
rect 316 411 325 1153
rect 334 510 343 1444
rect 352 1300 361 1746
rect 352 1295 356 1300
rect 352 599 361 1295
rect 370 1300 379 1935
rect 405 1431 837 1437
rect 370 698 380 1300
rect 405 718 415 1431
rect 425 1334 558 1339
rect 425 738 435 1334
rect 810 1312 837 1318
rect 445 1192 558 1197
rect 445 758 455 1192
rect 810 1170 837 1176
rect 465 1050 558 1055
rect 465 778 475 1050
rect 810 1028 837 1034
rect 810 886 837 892
rect 465 768 1998 778
rect 445 748 1978 758
rect 425 728 1958 738
rect 405 708 1937 718
rect 370 691 443 698
rect 352 593 414 599
rect 1927 575 1937 708
rect 334 503 415 510
rect 316 405 405 411
rect 1948 392 1958 728
rect 1924 387 1958 392
rect 298 315 415 322
rect 280 217 405 223
rect 1968 204 1978 748
rect 1938 199 1978 204
rect 262 127 408 133
rect 244 56 425 62
rect 1988 43 1998 768
rect 1918 38 1998 43
rect 368 19 382 24
rect 390 19 405 24
<< m2contact >>
rect 320 1153 325 1158
rect 280 764 289 771
rect 243 273 253 280
rect 356 1295 361 1300
rect 530 1295 535 1300
rect 530 1153 535 1158
rect 530 1011 537 1016
rect 530 908 539 913
rect 529 869 539 874
rect 382 19 390 24
<< metal2 >>
rect 361 1295 530 1300
rect 325 1153 530 1158
rect 280 1011 530 1016
rect 280 771 289 1011
rect 280 763 289 764
rect 308 908 530 913
rect 308 280 315 908
rect 382 869 529 874
rect 253 273 316 280
rect 382 24 390 869
use png  png_0
timestamp 1619529522
transform 0 -1 187 1 0 108
box -108 -66 1834 187
use sumblock  sumblock_0
timestamp 1619529573
transform 1 0 530 0 1 1249
box 0 -426 307 128
use carrygen  carrygen_0
timestamp 1619529550
transform 1 0 408 0 1 -5
box -26 0 1530 703
<< end >>
