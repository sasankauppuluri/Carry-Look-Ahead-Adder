magic
tech scmos
timestamp 1619529550
<< metal1 >>
rect -26 696 1351 703
rect -1 671 810 680
rect -1 604 6 671
rect 203 604 210 671
rect 324 659 447 665
rect 376 622 438 627
rect -26 598 33 604
rect 0 515 7 566
rect 174 531 180 601
rect 203 598 237 604
rect 376 596 383 622
rect 599 604 605 671
rect 724 659 789 665
rect 804 604 810 671
rect 928 659 1029 665
rect 1103 659 1199 665
rect 1147 622 1187 627
rect 1345 622 1351 696
rect 599 598 637 604
rect 804 598 842 604
rect 376 575 436 580
rect 214 537 252 542
rect 376 531 383 575
rect 174 525 383 531
rect 567 534 572 585
rect 981 580 988 601
rect 1147 580 1154 622
rect 1315 580 1321 585
rect 1458 580 1529 585
rect 981 575 1018 580
rect 588 537 657 542
rect 728 537 862 542
rect 933 537 1032 542
rect 1162 534 1169 580
rect 1315 575 1352 580
rect 1268 537 1367 542
rect 567 529 1169 534
rect -26 508 816 515
rect -2 483 605 492
rect -2 416 5 483
rect 121 471 190 477
rect 203 416 210 483
rect 324 471 461 477
rect 376 434 438 439
rect -26 410 33 416
rect 203 410 237 416
rect 376 408 383 434
rect 599 416 605 483
rect 719 471 789 477
rect 810 434 816 508
rect 902 471 1003 477
rect 947 434 993 439
rect 599 410 637 416
rect 0 327 7 378
rect 174 342 180 408
rect 376 387 436 392
rect 227 349 257 354
rect 376 342 383 387
rect 174 337 383 342
rect 567 346 572 397
rect 777 393 783 408
rect 777 387 817 393
rect 947 392 953 434
rect 1097 392 1530 397
rect 625 349 657 354
rect 728 349 831 354
rect 968 346 973 392
rect 567 341 973 346
rect -26 320 605 327
rect -2 295 210 304
rect -2 228 5 295
rect 121 283 189 289
rect 203 228 210 295
rect 323 283 447 289
rect 376 246 438 251
rect 599 246 605 320
rect -26 222 39 228
rect 203 222 238 228
rect 376 220 383 246
rect 0 138 7 190
rect 174 157 180 220
rect 567 204 572 209
rect 711 204 1530 209
rect 376 199 436 204
rect 567 199 606 204
rect 227 161 252 166
rect 376 157 383 199
rect 520 161 620 166
rect 174 152 383 157
rect -26 132 227 138
rect 121 122 210 128
rect 222 85 227 132
rect -26 61 34 67
rect 174 43 180 59
rect 330 43 1530 48
rect 174 38 210 43
rect -26 24 33 29
rect 125 0 243 5
<< m2contact >>
rect 39 659 46 665
rect 119 659 126 665
rect 242 659 249 665
rect 520 659 526 665
rect 125 537 132 543
rect 642 659 648 665
rect 789 659 795 665
rect 847 659 853 665
rect 1270 659 1275 665
rect 1358 659 1363 665
rect 777 596 783 601
rect 207 537 214 543
rect 328 537 335 542
rect 445 537 452 542
rect 519 537 524 542
rect 583 537 588 542
rect 1100 537 1106 542
rect 1460 557 1465 562
rect 1194 537 1200 542
rect 39 471 46 477
rect 190 471 196 477
rect 242 471 248 477
rect 519 471 526 477
rect 174 408 180 413
rect 642 471 649 477
rect 789 471 795 477
rect 823 471 829 477
rect 777 408 783 413
rect 125 349 132 355
rect 220 349 227 355
rect 328 349 335 354
rect 445 349 452 354
rect 517 349 524 354
rect 618 349 625 354
rect 900 349 905 354
rect 1099 369 1104 374
rect 1000 349 1005 354
rect 39 283 46 289
rect 189 283 195 289
rect 242 283 248 289
rect 521 283 526 289
rect 612 283 617 289
rect 174 220 180 225
rect 125 161 132 166
rect 220 161 227 166
rect 328 161 335 166
rect 714 181 719 186
rect 445 161 450 166
rect 39 122 46 128
rect 210 122 216 128
rect 235 122 241 128
rect 174 59 180 64
rect 337 20 342 25
<< metal2 >>
rect 777 684 1023 691
rect 15 659 39 665
rect 126 659 242 665
rect 526 659 642 665
rect 15 477 22 659
rect 777 601 783 684
rect 795 659 847 665
rect 1020 622 1023 684
rect 1275 659 1358 665
rect 132 537 207 543
rect 236 523 243 566
rect 335 537 445 542
rect 524 537 583 542
rect 636 526 643 566
rect 841 526 848 566
rect 1106 537 1194 542
rect 174 519 243 523
rect 15 471 39 477
rect 15 289 22 471
rect 174 413 180 519
rect 438 518 643 526
rect 777 518 848 526
rect 196 471 242 477
rect 438 434 441 518
rect 526 471 642 477
rect 777 413 783 518
rect 795 471 823 477
rect 132 349 220 355
rect 236 335 243 378
rect 335 349 445 354
rect 524 349 618 354
rect 636 338 643 378
rect 1460 374 1465 557
rect 1104 369 1465 374
rect 905 349 1000 354
rect 174 331 243 335
rect 15 283 39 289
rect 15 128 22 283
rect 174 225 180 331
rect 438 330 643 338
rect 195 283 242 289
rect 438 246 441 330
rect 526 283 612 289
rect 132 161 220 166
rect 236 151 243 190
rect 1099 186 1104 369
rect 719 181 1104 186
rect 335 161 445 166
rect 174 147 243 151
rect 15 122 39 128
rect 174 64 180 147
rect 216 122 235 128
rect 714 24 719 181
rect 342 20 719 24
use andgate  andgate_6
timestamp 1618893190
transform 1 0 115 0 1 573
box -115 -36 65 92
use andgate  andgate_7
timestamp 1618893190
transform 1 0 318 0 1 573
box -115 -36 65 92
use orgate  orgate_6
timestamp 1618893311
transform 1 0 516 0 1 557
box -103 -20 56 108
use andgate  andgate_8
timestamp 1618893190
transform 1 0 718 0 1 573
box -115 -36 65 92
use andgate  andgate_9
timestamp 1618893190
transform 1 0 923 0 1 573
box -115 -36 65 92
use orgate  orgate_7
timestamp 1618893311
transform 1 0 1098 0 1 557
box -103 -20 56 108
use orgate  orgate_8
timestamp 1618893311
transform 1 0 1265 0 1 557
box -103 -20 56 108
use orgate  orgate_9
timestamp 1618893311
transform 1 0 1432 0 1 557
box -103 -20 56 108
use andgate  andgate_3
timestamp 1618893190
transform 1 0 115 0 1 385
box -115 -36 65 92
use andgate  andgate_4
timestamp 1618893190
transform 1 0 318 0 1 385
box -115 -36 65 92
use orgate  orgate_3
timestamp 1618893311
transform 1 0 516 0 1 369
box -103 -20 56 108
use andgate  andgate_5
timestamp 1618893190
transform 1 0 718 0 1 385
box -115 -36 65 92
use orgate  orgate_4
timestamp 1618893311
transform 1 0 897 0 1 369
box -103 -20 56 108
use orgate  orgate_5
timestamp 1618893311
transform 1 0 1071 0 1 369
box -103 -20 56 108
use andgate  andgate_1
timestamp 1618893190
transform 1 0 115 0 1 197
box -115 -36 65 92
use andgate  andgate_2
timestamp 1618893190
transform 1 0 318 0 1 197
box -115 -36 65 92
use orgate  orgate_1
timestamp 1618893311
transform 1 0 516 0 1 181
box -103 -20 56 108
use orgate  orgate_2
timestamp 1618893311
transform 1 0 686 0 1 181
box -103 -20 56 108
use andgate  andgate_0
timestamp 1618893190
transform 1 0 115 0 1 36
box -115 -36 65 92
use orgate  orgate_0
timestamp 1618893311
transform 1 0 309 0 1 20
box -103 -20 56 108
<< end >>
