magic
tech scmos
timestamp 1618846832
<< nwell >>
rect -71 38 -43 70
rect -37 30 -9 62
rect 41 38 69 70
rect 75 30 103 62
<< ntransistor >>
rect -58 -20 -56 -10
rect -24 -12 -22 -2
rect 54 -20 56 -10
rect 88 -12 90 -2
<< ptransistor >>
rect -58 44 -56 64
rect -24 36 -22 56
rect 54 44 56 64
rect 88 36 90 56
<< ndiffusion >>
rect -59 -20 -58 -10
rect -56 -20 -55 -10
rect -25 -12 -24 -2
rect -22 -12 -21 -2
rect 53 -20 54 -10
rect 56 -20 57 -10
rect 87 -12 88 -2
rect 90 -12 91 -2
<< pdiffusion >>
rect -59 44 -58 64
rect -56 44 -55 64
rect -25 36 -24 56
rect -22 36 -21 56
rect 53 44 54 64
rect 56 44 57 64
rect 87 36 88 56
rect 90 36 91 56
<< ndcontact >>
rect -64 -20 -59 -10
rect -55 -20 -50 -10
rect -30 -12 -25 -2
rect -21 -12 -16 -2
rect 48 -20 53 -10
rect 57 -20 62 -10
rect 82 -12 87 -2
rect 91 -12 96 -2
<< pdcontact >>
rect -64 44 -59 64
rect -55 44 -50 64
rect -30 36 -25 56
rect -21 36 -16 56
rect 48 44 53 64
rect 57 44 62 64
rect 82 36 87 56
rect 91 36 96 56
<< polysilicon >>
rect -58 64 -56 67
rect 54 64 56 67
rect -24 56 -22 59
rect -58 30 -56 44
rect 88 56 90 59
rect -24 21 -22 36
rect 54 30 56 44
rect 88 21 90 36
rect -24 -2 -22 6
rect 88 -2 90 6
rect -58 -10 -56 -2
rect 54 -10 56 -2
rect -24 -16 -22 -12
rect 88 -16 90 -12
rect -58 -24 -56 -20
rect 54 -24 56 -20
<< polycontact >>
rect -64 32 -58 37
rect -30 23 -24 28
rect 48 32 54 37
rect 82 23 88 28
rect -30 1 -24 6
rect 82 1 88 6
rect -64 -7 -58 -2
rect 48 -7 54 -2
<< metal1 >>
rect -106 69 69 75
rect -64 64 -59 69
rect 5 64 9 69
rect 48 64 53 69
rect -50 44 -30 51
rect -77 37 -72 42
rect -130 32 -111 37
rect -90 32 -64 37
rect 62 44 82 51
rect -119 6 -114 32
rect -37 23 -30 28
rect -21 16 -16 36
rect 46 32 48 37
rect 36 23 82 28
rect -106 13 -90 14
rect -85 13 -78 14
rect -119 1 -30 6
rect -21 -2 -16 10
rect -142 -7 -76 -2
rect -70 -7 -64 -2
rect -55 -10 -30 -6
rect -90 -48 -85 -17
rect -64 -48 -59 -20
rect 12 -48 17 2
rect 36 -2 39 23
rect 91 16 96 36
rect 96 10 138 16
rect 77 1 82 6
rect 91 -2 96 10
rect 36 -7 48 -2
rect 57 -10 82 -6
rect 48 -48 53 -20
rect -90 -53 69 -48
<< m2contact >>
rect -77 42 -72 47
rect -107 32 -102 37
rect -42 23 -37 28
rect 41 32 46 37
rect 0 23 5 28
rect -90 9 -85 14
rect -21 10 -16 16
rect -76 -7 -70 -2
rect -90 -17 -85 -12
rect 91 10 96 16
rect 70 1 77 6
<< metal2 >>
rect -72 42 113 47
rect -102 32 41 37
rect -76 23 -42 28
rect -37 23 0 28
rect -90 -12 -85 9
rect -76 -2 -70 23
rect -16 10 91 16
rect 107 6 113 42
rect 77 1 113 6
use inverter  inverter_1
timestamp 1618833239
transform 1 0 -93 0 1 45
box -18 -36 21 30
use inverter  inverter_0
timestamp 1618833239
transform 1 0 18 0 1 36
box -18 -36 21 30
<< end >>
