* SPICE3 file created from pngblock.ext - technology: scmos

.option scale=0.09u

M1000 m1_465_n34# andgate_0/a_n61_61# a_537_97# andgate_0/inverter_0/w_n13_n7# pfet w=20 l=2
+  ad=120 pd=52 as=3360 ps=1456
M1001 m1_465_n34# andgate_0/a_n61_61# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=1440 ps=768
M1002 andgate_0/a_n61_61# m1_11_142# a_537_97# andgate_0/w_n76_50# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1003 andgate_0/a_n61_61# m1_0_46# a_537_97# andgate_0/w_n42_50# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 andgate_0/a_n61_61# m1_11_142# andgate_0/a_n58_n26# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=120 ps=64
M1005 andgate_0/a_n58_n26# m1_0_46# a_537_72# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 xorgate_0/a_48_n7# m1_0_46# a_537_97# xorgate_0/inverter_0/w_n13_n7# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1007 xorgate_0/a_48_n7# m1_0_46# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1008 xorgate_0/a_n64_32# m1_11_142# a_537_97# xorgate_0/inverter_1/w_n13_n7# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1009 xorgate_0/a_n64_32# m1_11_142# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1010 xorgate_0/a_n56_44# xorgate_0/a_n64_32# a_537_97# xorgate_0/w_n71_38# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1011 m1_272_n34# m1_0_46# xorgate_0/a_n56_44# xorgate_0/w_n37_30# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1012 xorgate_0/a_56_44# m1_11_142# a_537_97# xorgate_0/w_41_38# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1013 m1_272_n34# xorgate_0/a_48_n7# xorgate_0/a_56_44# xorgate_0/w_75_30# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 xorgate_0/a_n56_n20# m1_0_46# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1015 m1_272_n34# m1_11_142# xorgate_0/a_n56_n20# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1016 xorgate_0/a_56_n20# xorgate_0/a_48_n7# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1017 m1_272_n34# xorgate_0/a_n64_32# xorgate_0/a_56_n20# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 a_545_72# a_537_85# a_537_97# w_530_91# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1019 a_580_97# a_545_72# a_537_97# w_565_91# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1020 a_614_41# a_572_46# a_580_97# w_599_83# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1021 a_545_72# a_537_85# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1022 a_656_63# a_572_46# a_537_97# w_641_82# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1023 a_692_97# a_537_85# a_537_97# w_677_91# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1024 a_614_41# a_656_63# a_692_97# w_711_83# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 a_841_97# a_537_85# a_537_97# w_826_86# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1026 a_841_97# a_572_46# a_537_97# w_860_86# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 a_1038_72# a_1030_85# a_537_97# w_1023_91# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1028 a_1073_97# a_1038_72# a_537_97# w_1058_91# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1029 a_656_63# a_572_46# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1030 a_922_46# a_841_97# a_537_97# w_907_65# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1031 a_1107_41# a_1065_46# a_1073_97# w_1092_83# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1032 a_1038_72# a_1030_85# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1033 a_1149_63# a_1065_46# a_537_97# w_1134_82# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1034 a_1185_97# a_1030_85# a_537_97# w_1170_91# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1035 a_1107_41# a_1149_63# a_1185_97# w_1204_83# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 a_1334_97# a_1030_85# a_537_97# w_1319_86# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1037 a_1334_97# a_1065_46# a_537_97# w_1353_86# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 a_1532_72# a_1524_85# a_537_97# w_1517_91# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1039 a_1567_97# a_1532_72# a_537_97# w_1552_91# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1040 a_1149_63# a_1065_46# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1041 a_1415_46# a_1334_97# a_537_97# w_1400_65# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1042 a_1601_41# a_1559_46# a_1567_97# w_1586_83# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1043 a_1532_72# a_1524_85# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1044 a_1643_63# a_1559_46# a_537_97# w_1628_82# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1045 a_1679_97# a_1524_85# a_537_97# w_1664_91# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1046 a_1601_41# a_1643_63# a_1679_97# w_1698_83# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 a_1828_97# a_1524_85# a_537_97# w_1813_86# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1048 a_1828_97# a_1559_46# a_537_97# w_1847_86# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 a_580_33# a_572_46# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1050 a_614_41# a_537_85# a_580_33# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1051 a_692_33# a_656_63# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1052 a_614_41# a_545_72# a_692_33# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 a_841_97# a_537_85# a_844_10# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=120 ps=64
M1054 a_922_46# a_841_97# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1055 a_1643_63# a_1559_46# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1056 a_1909_46# a_1828_97# a_537_97# w_1894_65# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1057 a_1073_33# a_1065_46# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1058 a_1107_41# a_1030_85# a_1073_33# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1059 a_1185_33# a_1149_63# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1060 a_1107_41# a_1038_72# a_1185_33# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 a_1334_97# a_1030_85# a_1337_10# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=120 ps=64
M1062 a_1415_46# a_1334_97# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1063 a_1567_33# a_1559_46# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1064 a_1601_41# a_1524_85# a_1567_33# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1065 a_1679_33# a_1643_63# a_537_72# Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1066 a_1601_41# a_1532_72# a_1679_33# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_1828_97# a_1524_85# a_1831_10# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=120 ps=64
M1068 a_1909_46# a_1828_97# a_537_72# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1069 a_844_10# a_572_46# a_537_72# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 a_1337_10# a_1065_46# a_537_72# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 a_1831_10# a_1559_46# a_537_72# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_1073_97# w_1092_83# 0.1fF
C1 a_537_85# w_641_82# 0.2fF
C2 a_1831_10# a_537_72# 0.1fF
C3 a_1532_72# a_1524_85# 0.5fF
C4 a_841_97# w_826_86# 0.1fF
C5 a_1415_46# w_1400_65# 0.0fF
C6 m1_0_46# andgate_0/w_n42_50# 0.1fF
C7 a_922_46# a_537_72# 0.3fF
C8 a_1038_72# w_1204_83# 0.1fF
C9 a_1334_97# w_1353_86# 0.1fF
C10 a_1065_46# w_1353_86# 0.1fF
C11 w_1664_91# a_537_97# 0.1fF
C12 a_1185_97# a_537_97# 0.2fF
C13 a_1149_63# a_537_97# 0.2fF
C14 xorgate_0/a_56_n20# xorgate_0/a_n64_32# 0.1fF
C15 w_907_65# a_537_97# 0.1fF
C16 xorgate_0/a_n56_44# a_537_97# 0.2fF
C17 xorgate_0/a_n64_32# xorgate_0/a_48_n7# 0.0fF
C18 m1_465_n34# a_537_97# 0.2fF
C19 a_537_85# a_537_72# 0.6fF
C20 a_1601_41# a_537_72# 0.2fF
C21 m1_11_142# xorgate_0/inverter_0/w_n13_n7# 0.0fF
C22 m1_0_46# a_537_72# 0.4fF
C23 a_692_33# a_614_41# 0.1fF
C24 a_580_33# a_614_41# 0.1fF
C25 a_1679_97# a_1532_72# 0.4fF
C26 a_1038_72# w_1134_82# 0.2fF
C27 a_1038_72# w_1058_91# 0.2fF
C28 a_614_41# a_545_72# 0.6fF
C29 a_922_46# w_907_65# 0.0fF
C30 a_545_72# w_677_91# 0.2fF
C31 a_922_46# a_537_97# 0.2fF
C32 m1_272_n34# xorgate_0/a_n64_32# 0.6fF
C33 andgate_0/w_n76_50# a_537_97# 0.1fF
C34 a_692_33# a_545_72# 0.1fF
C35 m1_272_n34# xorgate_0/w_n37_30# 0.0fF
C36 a_1679_33# a_1601_41# 0.1fF
C37 a_1337_10# a_1065_46# 0.2fF
C38 a_1337_10# a_1334_97# 0.1fF
C39 a_1185_33# a_1038_72# 0.1fF
C40 a_1337_10# a_1030_85# 0.1fF
C41 a_1567_33# a_1559_46# 0.0fF
C42 a_656_63# a_572_46# 0.1fF
C43 a_1107_41# a_1065_46# 0.2fF
C44 a_1107_41# a_1030_85# 0.2fF
C45 a_1073_97# a_1038_72# 0.4fF
C46 a_1601_41# w_1698_83# 0.0fF
C47 a_537_85# a_537_97# 0.5fF
C48 w_860_86# a_537_97# 0.1fF
C49 xorgate_0/a_56_44# a_537_97# 0.2fF
C50 m1_0_46# a_537_97# 0.2fF
C51 andgate_0/a_n58_n26# m1_11_142# 0.1fF
C52 a_1532_72# w_1552_91# 0.2fF
C53 a_1073_97# w_1058_91# 0.1fF
C54 a_841_97# a_572_46# 0.3fF
C55 a_1601_41# w_1586_83# 0.0fF
C56 xorgate_0/a_56_44# xorgate_0/w_75_30# 0.1fF
C57 a_1567_33# a_1524_85# 0.2fF
C58 a_614_41# a_692_97# 0.2fF
C59 a_1334_97# a_537_72# 0.1fF
C60 a_1065_46# a_537_72# 0.4fF
C61 a_1030_85# a_537_72# 0.6fF
C62 a_692_97# w_677_91# 0.1fF
C63 a_1567_97# a_537_97# 0.2fF
C64 a_1828_97# a_537_72# 0.1fF
C65 w_1847_86# a_537_97# 0.1fF
C66 w_826_86# a_537_97# 0.1fF
C67 xorgate_0/a_56_n20# a_537_72# 0.1fF
C68 xorgate_0/a_n56_n20# a_537_72# 0.1fF
C69 xorgate_0/a_n64_32# xorgate_0/inverter_0/w_n13_n7# 0.0fF
C70 xorgate_0/a_48_n7# a_537_72# 0.2fF
C71 a_1643_63# w_1628_82# 0.0fF
C72 a_1559_46# w_1628_82# 0.1fF
C73 a_1107_41# w_1092_83# 0.0fF
C74 a_572_46# w_641_82# 0.1fF
C75 a_1524_85# w_1517_91# 0.1fF
C76 a_1567_97# w_1586_83# 0.1fF
C77 a_692_97# a_545_72# 0.4fF
C78 a_1415_46# a_537_72# 0.3fF
C79 xorgate_0/w_41_38# m1_11_142# 0.1fF
C80 m1_272_n34# a_537_72# 0.2fF
C81 a_1149_63# a_1065_46# 0.1fF
C82 a_1149_63# a_1030_85# 0.2fF
C83 a_656_63# a_614_41# 0.3fF
C84 a_1601_41# a_1567_97# 0.2fF
C85 w_1813_86# a_537_97# 0.1fF
C86 a_1828_97# a_537_97# 0.6fF
C87 a_1334_97# a_537_97# 0.6fF
C88 a_1065_46# a_537_97# 0.4fF
C89 a_1030_85# a_537_97# 0.5fF
C90 w_565_91# a_537_97# 0.1fF
C91 a_1524_85# w_1628_82# 0.2fF
C92 xorgate_0/a_48_n7# a_537_97# 0.2fF
C93 andgate_0/a_n58_n26# andgate_0/a_n61_61# 0.1fF
C94 a_572_46# a_537_72# 0.4fF
C95 a_537_85# w_826_86# 0.1fF
C96 a_1643_63# a_537_72# 0.3fF
C97 a_1559_46# a_537_72# 0.4fF
C98 a_1831_10# a_1828_97# 0.1fF
C99 a_844_10# a_841_97# 0.1fF
C100 a_692_33# a_656_63# 0.0fF
C101 a_656_63# a_545_72# 0.1fF
C102 a_1415_46# a_537_97# 0.2fF
C103 a_545_72# w_530_91# 0.0fF
C104 w_1894_65# a_537_97# 0.1fF
C105 xorgate_0/a_n56_44# m1_272_n34# 0.2fF
C106 xorgate_0/w_75_30# xorgate_0/a_48_n7# 0.1fF
C107 a_1524_85# a_537_72# 0.6fF
C108 a_1532_72# w_1517_91# 0.0fF
C109 m1_272_n34# xorgate_0/w_75_30# 0.0fF
C110 a_1679_33# a_1643_63# 0.0fF
C111 a_1643_63# w_1698_83# 0.1fF
C112 a_1185_97# w_1170_91# 0.1fF
C113 a_1107_41# w_1204_83# 0.0fF
C114 a_1107_41# a_1038_72# 0.6fF
C115 a_1643_63# a_537_97# 0.2fF
C116 a_1559_46# a_537_97# 0.4fF
C117 a_580_97# a_537_97# 0.2fF
C118 a_572_46# a_537_97# 0.4fF
C119 w_1170_91# a_537_97# 0.1fF
C120 xorgate_0/w_41_38# xorgate_0/a_n64_32# 0.2fF
C121 xorgate_0/a_n56_n20# m1_0_46# 0.0fF
C122 xorgate_0/a_n64_32# m1_11_142# 0.5fF
C123 xorgate_0/a_48_n7# m1_0_46# 0.1fF
C124 m1_11_142# andgate_0/a_n61_61# 0.1fF
C125 a_1831_10# a_1559_46# 0.2fF
C126 a_1559_46# w_1586_83# 0.1fF
C127 a_537_85# w_599_83# 0.2fF
C128 a_1532_72# w_1628_82# 0.2fF
C129 a_545_72# w_641_82# 0.2fF
C130 xorgate_0/w_n37_30# m1_11_142# 0.2fF
C131 xorgate_0/a_56_44# m1_272_n34# 0.2fF
C132 m1_272_n34# m1_0_46# 0.2fF
C133 m1_11_142# xorgate_0/inverter_1/w_n13_n7# 0.1fF
C134 a_1828_97# w_1847_86# 0.1fF
C135 a_844_10# a_537_72# 0.1fF
C136 a_1524_85# w_1664_91# 0.1fF
C137 a_614_41# a_537_72# 0.2fF
C138 a_1909_46# a_537_72# 0.1fF
C139 a_1038_72# a_537_72# 0.1fF
C140 a_1524_85# a_537_97# 0.5fF
C141 w_1023_91# a_537_97# 0.1fF
C142 xorgate_0/w_n71_38# xorgate_0/a_n64_32# 0.2fF
C143 xorgate_0/inverter_0/w_n13_n7# a_537_97# 0.1fF
C144 andgate_0/a_n58_n26# a_537_72# 0.1fF
C145 a_1185_33# a_1107_41# 0.1fF
C146 a_1643_63# a_1601_41# 0.3fF
C147 a_580_97# a_537_85# 0.1fF
C148 a_572_46# a_537_85# 2.5fF
C149 a_1601_41# a_1559_46# 0.2fF
C150 a_1107_41# a_1073_97# 0.2fF
C151 a_1831_10# a_1524_85# 0.1fF
C152 a_572_46# w_860_86# 0.1fF
C153 a_692_33# a_537_72# 0.1fF
C154 a_580_33# a_537_72# 0.1fF
C155 a_1524_85# w_1586_83# 0.2fF
C156 a_1532_72# a_537_72# 0.1fF
C157 a_545_72# a_537_72# 0.1fF
C158 a_1334_97# a_1065_46# 0.3fF
C159 a_1334_97# a_1030_85# 0.1fF
C160 a_1065_46# a_1030_85# 2.5fF
C161 a_1185_97# w_1204_83# 0.1fF
C162 a_1149_63# w_1204_83# 0.1fF
C163 a_1828_97# w_1813_86# 0.1fF
C164 a_1185_97# a_1038_72# 0.4fF
C165 a_1679_97# w_1698_83# 0.1fF
C166 a_1679_97# w_1664_91# 0.1fF
C167 a_1149_63# a_1038_72# 0.1fF
C168 a_1679_97# a_537_97# 0.2fF
C169 a_1909_46# a_537_97# 0.2fF
C170 a_1038_72# a_537_97# 0.6fF
C171 a_1073_33# a_1107_41# 0.1fF
C172 a_1601_41# a_1524_85# 0.2fF
C173 a_614_41# w_711_83# 0.0fF
C174 a_1559_46# w_1847_86# 0.1fF
C175 w_1319_86# a_537_97# 0.1fF
C176 w_677_91# a_537_97# 0.1fF
C177 a_1185_33# a_537_72# 0.1fF
C178 xorgate_0/a_56_n20# xorgate_0/a_48_n7# 0.0fF
C179 m1_11_142# a_537_72# 0.4fF
C180 xorgate_0/inverter_0/w_n13_n7# m1_0_46# 0.1fF
C181 a_1828_97# w_1894_65# 0.1fF
C182 a_1334_97# a_1415_46# 0.1fF
C183 a_1679_33# a_1532_72# 0.1fF
C184 a_1149_63# w_1134_82# 0.0fF
C185 a_1532_72# w_1698_83# 0.1fF
C186 a_1532_72# w_1664_91# 0.2fF
C187 a_545_72# a_537_97# 0.6fF
C188 a_1532_72# a_537_97# 0.6fF
C189 w_1134_82# a_537_97# 0.1fF
C190 w_1058_91# a_537_97# 0.1fF
C191 a_545_72# w_711_83# 0.1fF
C192 xorgate_0/w_n37_30# xorgate_0/a_n64_32# 0.1fF
C193 xorgate_0/a_56_n20# m1_272_n34# 0.1fF
C194 xorgate_0/a_n56_n20# m1_272_n34# 0.1fF
C195 m1_272_n34# xorgate_0/a_48_n7# 0.2fF
C196 xorgate_0/a_n64_32# xorgate_0/inverter_1/w_n13_n7# 0.0fF
C197 a_1567_97# a_1524_85# 0.1fF
C198 a_1073_33# a_537_72# 0.1fF
C199 a_1532_72# w_1586_83# 0.1fF
C200 a_1828_97# a_1559_46# 0.3fF
C201 a_1679_97# a_1601_41# 0.2fF
C202 a_844_10# a_537_85# 0.1fF
C203 a_1185_33# a_1149_63# 0.0fF
C204 a_580_97# w_565_91# 0.1fF
C205 a_1030_85# w_1170_91# 0.1fF
C206 a_1065_46# w_1092_83# 0.1fF
C207 a_614_41# a_537_85# 0.2fF
C208 a_1030_85# w_1092_83# 0.2fF
C209 a_1073_97# a_537_97# 0.2fF
C210 a_656_63# w_641_82# 0.0fF
C211 a_537_85# w_677_91# 0.1fF
C212 w_1552_91# a_537_97# 0.1fF
C213 xorgate_0/a_n56_44# m1_11_142# 0.1fF
C214 xorgate_0/w_41_38# a_537_97# 0.1fF
C215 m1_11_142# a_537_97# 0.2fF
C216 andgate_0/a_n61_61# andgate_0/w_n42_50# 0.1fF
C217 andgate_0/a_n58_n26# m1_0_46# 0.2fF
C218 andgate_0/a_n61_61# andgate_0/inverter_0/w_n13_n7# 0.1fF
C219 a_1601_41# a_1532_72# 0.6fF
C220 a_580_33# a_537_85# 0.2fF
C221 a_580_97# w_599_83# 0.1fF
C222 a_545_72# a_537_85# 0.5fF
C223 a_572_46# w_599_83# 0.1fF
C224 m1_11_142# andgate_0/w_n76_50# 0.1fF
C225 a_1828_97# a_1524_85# 0.1fF
C226 a_1524_85# w_1813_86# 0.1fF
C227 a_1567_33# a_537_72# 0.1fF
C228 a_692_97# w_711_83# 0.1fF
C229 a_1030_85# w_1023_91# 0.1fF
C230 w_1400_65# a_537_97# 0.1fF
C231 a_692_97# a_537_97# 0.2fF
C232 a_656_63# a_537_72# 0.3fF
C233 xorgate_0/a_n56_44# xorgate_0/w_n71_38# 0.1fF
C234 xorgate_0/w_n71_38# a_537_97# 0.1fF
C235 xorgate_0/a_n64_32# a_537_72# 0.1fF
C236 xorgate_0/inverter_0/w_n13_n7# xorgate_0/a_48_n7# 0.0fF
C237 andgate_0/a_n61_61# a_537_72# 0.1fF
C238 a_1643_63# a_1559_46# 0.1fF
C239 a_1567_97# a_1532_72# 0.4fF
C240 xorgate_0/a_56_44# xorgate_0/w_41_38# 0.1fF
C241 m1_11_142# m1_0_46# 2.3fF
C242 a_841_97# a_537_72# 0.1fF
C243 a_1909_46# a_1828_97# 0.1fF
C244 a_1334_97# w_1319_86# 0.1fF
C245 a_1030_85# w_1319_86# 0.1fF
C246 a_1065_46# a_1038_72# 0.0fF
C247 a_1030_85# a_1038_72# 0.5fF
C248 a_656_63# w_711_83# 0.1fF
C249 a_656_63# a_537_97# 0.2fF
C250 a_1643_63# a_1524_85# 0.2fF
C251 a_1559_46# a_1524_85# 2.5fF
C252 a_1567_97# w_1552_91# 0.1fF
C253 w_1353_86# a_537_97# 0.1fF
C254 a_1337_10# a_537_72# 0.1fF
C255 w_530_91# a_537_97# 0.1fF
C256 xorgate_0/a_n56_44# xorgate_0/a_n64_32# 0.4fF
C257 xorgate_0/a_n64_32# a_537_97# 0.5fF
C258 andgate_0/a_n61_61# a_537_97# 0.6fF
C259 m1_465_n34# andgate_0/a_n61_61# 0.1fF
C260 a_1107_41# a_537_72# 0.2fF
C261 a_1909_46# w_1894_65# 0.0fF
C262 a_614_41# w_599_83# 0.0fF
C263 a_1065_46# w_1134_82# 0.1fF
C264 a_1030_85# w_1134_82# 0.2fF
C265 a_841_97# w_907_65# 0.1fF
C266 a_545_72# w_565_91# 0.2fF
C267 a_841_97# a_537_97# 0.6fF
C268 w_1517_91# a_537_97# 0.1fF
C269 xorgate_0/a_n56_44# xorgate_0/w_n37_30# 0.1fF
C270 xorgate_0/w_75_30# xorgate_0/a_n64_32# 0.1fF
C271 xorgate_0/inverter_1/w_n13_n7# a_537_97# 0.1fF
C272 andgate_0/a_n61_61# andgate_0/w_n76_50# 0.1fF
C273 a_922_46# a_841_97# 0.1fF
C274 a_545_72# w_599_83# 0.1fF
C275 a_1149_63# a_1107_41# 0.3fF
C276 a_1567_33# a_1601_41# 0.1fF
C277 a_844_10# a_572_46# 0.2fF
C278 a_1038_72# w_1170_91# 0.2fF
C279 a_1073_97# a_1030_85# 0.1fF
C280 a_614_41# a_580_97# 0.2fF
C281 a_614_41# a_572_46# 0.2fF
C282 a_656_63# a_537_85# 0.2fF
C283 a_1185_97# a_1107_41# 0.2fF
C284 a_537_85# w_530_91# 0.1fF
C285 w_1628_82# a_537_97# 0.1fF
C286 a_1038_72# w_1092_83# 0.1fF
C287 xorgate_0/a_n56_n20# m1_11_142# 0.2fF
C288 w_641_82# a_537_97# 0.1fF
C289 xorgate_0/a_56_44# xorgate_0/a_n64_32# 0.4fF
C290 m1_11_142# xorgate_0/a_48_n7# 0.1fF
C291 xorgate_0/a_n64_32# m1_0_46# 0.0fF
C292 m1_0_46# andgate_0/a_n61_61# 0.3fF
C293 andgate_0/w_n42_50# a_537_97# 0.1fF
C294 m1_465_n34# andgate_0/inverter_0/w_n13_n7# 0.0fF
C295 a_537_97# andgate_0/inverter_0/w_n13_n7# 0.1fF
C296 a_1643_63# a_1532_72# 0.1fF
C297 a_580_33# a_572_46# 0.0fF
C298 a_841_97# a_537_85# 0.1fF
C299 a_580_97# a_545_72# 0.4fF
C300 a_572_46# a_545_72# 0.0fF
C301 a_841_97# w_860_86# 0.1fF
C302 a_1559_46# a_1532_72# 0.0fF
C303 m1_272_n34# m1_11_142# 0.2fF
C304 xorgate_0/w_n37_30# m1_0_46# 0.1fF
C305 a_1073_33# a_1065_46# 0.0fF
C306 a_1073_33# a_1030_85# 0.2fF
C307 a_1038_72# w_1023_91# 0.0fF
C308 a_1334_97# w_1400_65# 0.1fF
C309 a_1679_33# a_537_72# 0.1fF
C310 a_1149_63# a_537_72# 0.3fF
C311 m1_465_n34# a_537_72# 0.3fF
C312 a_1831_10# gnd! 0.1fF
C313 a_1679_33# gnd! 0.1fF
C314 a_1567_33# gnd! 0.1fF
C315 a_1337_10# gnd! 0.1fF
C316 a_1185_33# gnd! 0.1fF
C317 a_1073_33# gnd! 0.1fF
C318 a_1909_46# gnd! 0.6fF
C319 a_844_10# gnd! 0.1fF
C320 a_692_33# gnd! 0.1fF
C321 a_580_33# gnd! 0.1fF
C322 a_1828_97# gnd! 0.6fF
C323 a_1679_97# gnd! 0.0fF
C324 a_1643_63# gnd! 0.6fF
C325 a_1601_41# gnd! 1.9fF
C326 a_1415_46# gnd! 0.6fF
C327 a_1567_97# gnd! 0.0fF
C328 a_1334_97# gnd! 0.6fF
C329 a_1185_97# gnd! 0.0fF
C330 a_1149_63# gnd! 0.6fF
C331 a_1107_41# gnd! 1.9fF
C332 a_922_46# gnd! 0.6fF
C333 a_1073_97# gnd! 0.0fF
C334 a_841_97# gnd! 0.6fF
C335 a_692_97# gnd! 0.0fF
C336 a_656_63# gnd! 0.6fF
C337 a_614_41# gnd! 1.9fF
C338 a_580_97# gnd! 0.0fF
C339 a_1559_46# gnd! 8.5fF
C340 a_1532_72# gnd! 1.7fF
C341 a_1524_85# gnd! 6.9fF
C342 a_1065_46# gnd! 8.5fF
C343 a_1038_72# gnd! 1.7fF
C344 a_1030_85# gnd! 6.9fF
C345 a_572_46# gnd! 8.5fF
C346 a_545_72# gnd! 1.7fF
C347 a_537_85# gnd! 6.9fF
C348 w_1894_65# gnd! 0.9fF
C349 w_1847_86# gnd! 1.0fF
C350 w_1813_86# gnd! 1.0fF
C351 w_1698_83# gnd! 0.9fF
C352 w_1664_91# gnd! 0.9fF
C353 w_1628_82# gnd! 0.9fF
C354 w_1586_83# gnd! 0.9fF
C355 w_1552_91# gnd! 0.9fF
C356 w_1517_91# gnd! 0.9fF
C357 w_1400_65# gnd! 0.9fF
C358 w_1353_86# gnd! 1.0fF
C359 w_1319_86# gnd! 1.0fF
C360 w_1204_83# gnd! 0.9fF
C361 w_1170_91# gnd! 0.9fF
C362 w_1134_82# gnd! 0.9fF
C363 w_1092_83# gnd! 0.9fF
C364 w_1058_91# gnd! 0.9fF
C365 w_1023_91# gnd! 0.9fF
C366 w_907_65# gnd! 0.9fF
C367 w_860_86# gnd! 1.0fF
C368 w_826_86# gnd! 1.0fF
C369 w_711_83# gnd! 0.9fF
C370 w_677_91# gnd! 0.9fF
C371 w_641_82# gnd! 0.9fF
C372 w_599_83# gnd! 0.9fF
C373 w_565_91# gnd! 0.9fF
C374 w_530_91# gnd! 0.9fF
C375 xorgate_0/a_56_n20# gnd! 0.1fF
C376 xorgate_0/a_n56_n20# gnd! 0.1fF
C377 xorgate_0/a_56_44# gnd! 0.0fF
C378 m1_272_n34# gnd! 2.1fF
C379 xorgate_0/a_n56_44# gnd! 0.0fF
C380 xorgate_0/w_75_30# gnd! 0.9fF
C381 xorgate_0/w_41_38# gnd! 0.9fF
C382 xorgate_0/w_n37_30# gnd! 0.9fF
C383 xorgate_0/w_n71_38# gnd! 0.9fF
C384 xorgate_0/a_n64_32# gnd! 1.0fF
C385 m1_11_142# gnd! 6.6fF
C386 xorgate_0/inverter_1/w_n13_n7# gnd! 0.9fF
C387 xorgate_0/a_48_n7# gnd! 0.6fF
C388 xorgate_0/inverter_0/w_n13_n7# gnd! 0.9fF
C389 andgate_0/a_n58_n26# gnd! 0.1fF
C390 m1_0_46# gnd! 7.8fF
C391 andgate_0/w_n42_50# gnd! 1.0fF
C392 andgate_0/w_n76_50# gnd! 1.0fF
C393 a_537_72# gnd! 18.7fF
C394 m1_465_n34# gnd! 0.6fF
C395 a_537_97# gnd! 13.4fF
C396 andgate_0/a_n61_61# gnd! 0.6fF
C397 andgate_0/inverter_0/w_n13_n7# gnd! 0.9fF
