magic
tech scmos
timestamp 1618833239
<< nwell >>
rect -13 -7 15 25
<< ntransistor >>
rect 0 -26 2 -16
<< ptransistor >>
rect 0 -1 2 19
<< ndiffusion >>
rect -1 -26 0 -16
rect 2 -26 3 -16
<< pdiffusion >>
rect -1 -1 0 19
rect 2 -1 3 19
<< ndcontact >>
rect -6 -26 -1 -16
rect 3 -26 8 -16
<< pdcontact >>
rect -6 -1 -1 19
rect 3 -1 8 19
<< polysilicon >>
rect 0 19 2 22
rect 0 -16 2 -1
rect 0 -30 2 -26
<< polycontact >>
rect -6 -13 0 -8
<< metal1 >>
rect -13 24 15 30
rect -6 19 -1 24
rect 3 -8 8 -1
rect -18 -13 -6 -8
rect 3 -13 21 -8
rect 3 -16 8 -13
rect -6 -32 -1 -26
rect -13 -36 15 -32
<< end >>
