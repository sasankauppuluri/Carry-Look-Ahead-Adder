magic
tech scmos
timestamp 1618855423
<< nwell >>
rect 530 91 558 123
rect 565 91 593 123
rect 599 83 627 115
rect 641 82 669 114
rect 677 91 705 123
rect 711 83 739 115
rect 826 86 854 123
rect 860 86 888 123
rect 907 65 935 97
rect 1023 91 1051 123
rect 1058 91 1086 123
rect 1092 83 1120 115
rect 1134 82 1162 114
rect 1170 91 1198 123
rect 1204 83 1232 115
rect 1319 86 1347 123
rect 1353 86 1381 123
rect 1400 65 1428 97
rect 1517 91 1545 123
rect 1552 91 1580 123
rect 1586 83 1614 115
rect 1628 82 1656 114
rect 1664 91 1692 123
rect 1698 83 1726 115
rect 1813 86 1841 123
rect 1847 86 1875 123
rect 1894 65 1922 97
<< ntransistor >>
rect 543 72 545 82
rect 654 63 656 73
rect 1036 72 1038 82
rect 1147 63 1149 73
rect 1530 72 1532 82
rect 578 33 580 43
rect 612 41 614 51
rect 690 33 692 43
rect 724 41 726 51
rect 851 41 853 51
rect 920 46 922 56
rect 1641 63 1643 73
rect 1071 33 1073 43
rect 1105 41 1107 51
rect 1183 33 1185 43
rect 1217 41 1219 51
rect 1344 41 1346 51
rect 1413 46 1415 56
rect 1565 33 1567 43
rect 1599 41 1601 51
rect 1677 33 1679 43
rect 1711 41 1713 51
rect 1838 41 1840 51
rect 1907 46 1909 56
rect 842 10 844 20
rect 1335 10 1337 20
rect 1829 10 1831 20
<< ptransistor >>
rect 543 97 545 117
rect 578 97 580 117
rect 612 89 614 109
rect 654 88 656 108
rect 690 97 692 117
rect 724 89 726 109
rect 839 97 841 117
rect 873 97 875 117
rect 1036 97 1038 117
rect 1071 97 1073 117
rect 920 71 922 91
rect 1105 89 1107 109
rect 1147 88 1149 108
rect 1183 97 1185 117
rect 1217 89 1219 109
rect 1332 97 1334 117
rect 1366 97 1368 117
rect 1530 97 1532 117
rect 1565 97 1567 117
rect 1413 71 1415 91
rect 1599 89 1601 109
rect 1641 88 1643 108
rect 1677 97 1679 117
rect 1711 89 1713 109
rect 1826 97 1828 117
rect 1860 97 1862 117
rect 1907 71 1909 91
<< ndiffusion >>
rect 542 72 543 82
rect 545 72 546 82
rect 653 63 654 73
rect 656 63 657 73
rect 1035 72 1036 82
rect 1038 72 1039 82
rect 1146 63 1147 73
rect 1149 63 1150 73
rect 1529 72 1530 82
rect 1532 72 1533 82
rect 577 33 578 43
rect 580 33 581 43
rect 611 41 612 51
rect 614 41 615 51
rect 689 33 690 43
rect 692 33 693 43
rect 723 41 724 51
rect 726 41 727 51
rect 850 41 851 51
rect 853 41 854 51
rect 919 46 920 56
rect 922 46 923 56
rect 1640 63 1641 73
rect 1643 63 1644 73
rect 1070 33 1071 43
rect 1073 33 1074 43
rect 1104 41 1105 51
rect 1107 41 1108 51
rect 1182 33 1183 43
rect 1185 33 1186 43
rect 1216 41 1217 51
rect 1219 41 1220 51
rect 1343 41 1344 51
rect 1346 41 1347 51
rect 1412 46 1413 56
rect 1415 46 1416 56
rect 1564 33 1565 43
rect 1567 33 1568 43
rect 1598 41 1599 51
rect 1601 41 1602 51
rect 1676 33 1677 43
rect 1679 33 1680 43
rect 1710 41 1711 51
rect 1713 41 1714 51
rect 1837 41 1838 51
rect 1840 41 1841 51
rect 1906 46 1907 56
rect 1909 46 1910 56
rect 841 10 842 20
rect 844 10 845 20
rect 1334 10 1335 20
rect 1337 10 1338 20
rect 1828 10 1829 20
rect 1831 10 1832 20
<< pdiffusion >>
rect 542 97 543 117
rect 545 97 546 117
rect 577 97 578 117
rect 580 97 581 117
rect 611 89 612 109
rect 614 89 615 109
rect 653 88 654 108
rect 656 88 657 108
rect 689 97 690 117
rect 692 97 693 117
rect 723 89 724 109
rect 726 89 727 109
rect 838 97 839 117
rect 841 97 842 117
rect 872 97 873 117
rect 875 97 876 117
rect 1035 97 1036 117
rect 1038 97 1039 117
rect 1070 97 1071 117
rect 1073 97 1074 117
rect 919 71 920 91
rect 922 71 923 91
rect 1104 89 1105 109
rect 1107 89 1108 109
rect 1146 88 1147 108
rect 1149 88 1150 108
rect 1182 97 1183 117
rect 1185 97 1186 117
rect 1216 89 1217 109
rect 1219 89 1220 109
rect 1331 97 1332 117
rect 1334 97 1335 117
rect 1365 97 1366 117
rect 1368 97 1369 117
rect 1529 97 1530 117
rect 1532 97 1533 117
rect 1564 97 1565 117
rect 1567 97 1568 117
rect 1412 71 1413 91
rect 1415 71 1416 91
rect 1598 89 1599 109
rect 1601 89 1602 109
rect 1640 88 1641 108
rect 1643 88 1644 108
rect 1676 97 1677 117
rect 1679 97 1680 117
rect 1710 89 1711 109
rect 1713 89 1714 109
rect 1825 97 1826 117
rect 1828 97 1829 117
rect 1859 97 1860 117
rect 1862 97 1863 117
rect 1906 71 1907 91
rect 1909 71 1910 91
<< ndcontact >>
rect 537 72 542 82
rect 546 72 551 82
rect 648 63 653 73
rect 657 63 662 73
rect 1030 72 1035 82
rect 1039 72 1044 82
rect 1141 63 1146 73
rect 1150 63 1155 73
rect 1524 72 1529 82
rect 1533 72 1538 82
rect 572 33 577 43
rect 581 33 586 43
rect 606 41 611 51
rect 615 41 620 51
rect 684 33 689 43
rect 693 33 698 43
rect 718 41 723 51
rect 727 41 732 51
rect 845 41 850 51
rect 854 41 859 51
rect 914 46 919 56
rect 923 46 928 56
rect 1635 63 1640 73
rect 1644 63 1649 73
rect 1065 33 1070 43
rect 1074 33 1079 43
rect 1099 41 1104 51
rect 1108 41 1113 51
rect 1177 33 1182 43
rect 1186 33 1191 43
rect 1211 41 1216 51
rect 1220 41 1225 51
rect 1338 41 1343 51
rect 1347 41 1352 51
rect 1407 46 1412 56
rect 1416 46 1421 56
rect 1559 33 1564 43
rect 1568 33 1573 43
rect 1593 41 1598 51
rect 1602 41 1607 51
rect 1671 33 1676 43
rect 1680 33 1685 43
rect 1705 41 1710 51
rect 1714 41 1719 51
rect 1832 41 1837 51
rect 1841 41 1846 51
rect 1901 46 1906 56
rect 1910 46 1915 56
rect 836 10 841 20
rect 845 10 850 20
rect 1329 10 1334 20
rect 1338 10 1343 20
rect 1823 10 1828 20
rect 1832 10 1837 20
<< pdcontact >>
rect 537 97 542 117
rect 546 97 551 117
rect 572 97 577 117
rect 581 97 586 117
rect 606 89 611 109
rect 615 89 620 109
rect 648 88 653 108
rect 657 88 662 108
rect 684 97 689 117
rect 693 97 698 117
rect 718 89 723 109
rect 727 89 732 109
rect 833 97 838 117
rect 842 97 847 117
rect 867 97 872 117
rect 876 97 881 117
rect 1030 97 1035 117
rect 1039 97 1044 117
rect 1065 97 1070 117
rect 1074 97 1079 117
rect 914 71 919 91
rect 923 71 928 91
rect 1099 89 1104 109
rect 1108 89 1113 109
rect 1141 88 1146 108
rect 1150 88 1155 108
rect 1177 97 1182 117
rect 1186 97 1191 117
rect 1211 89 1216 109
rect 1220 89 1225 109
rect 1326 97 1331 117
rect 1335 97 1340 117
rect 1360 97 1365 117
rect 1369 97 1374 117
rect 1524 97 1529 117
rect 1533 97 1538 117
rect 1559 97 1564 117
rect 1568 97 1573 117
rect 1407 71 1412 91
rect 1416 71 1421 91
rect 1593 89 1598 109
rect 1602 89 1607 109
rect 1635 88 1640 108
rect 1644 88 1649 108
rect 1671 97 1676 117
rect 1680 97 1685 117
rect 1705 89 1710 109
rect 1714 89 1719 109
rect 1820 97 1825 117
rect 1829 97 1834 117
rect 1854 97 1859 117
rect 1863 97 1868 117
rect 1901 71 1906 91
rect 1910 71 1915 91
<< polysilicon >>
rect 543 117 545 120
rect 578 117 580 120
rect 690 117 692 120
rect 839 117 841 120
rect 873 117 875 120
rect 1036 117 1038 120
rect 1071 117 1073 120
rect 1183 117 1185 120
rect 1332 117 1334 120
rect 1366 117 1368 120
rect 1530 117 1532 120
rect 1565 117 1567 120
rect 1677 117 1679 120
rect 1826 117 1828 120
rect 1860 117 1862 120
rect 612 109 614 112
rect 543 82 545 97
rect 578 83 580 97
rect 654 108 656 111
rect 612 74 614 89
rect 724 109 726 112
rect 654 73 656 88
rect 690 83 692 97
rect 1105 109 1107 112
rect 724 74 726 89
rect 839 76 841 97
rect 873 77 875 97
rect 920 91 922 94
rect 543 68 545 72
rect 1036 82 1038 97
rect 1071 83 1073 97
rect 1147 108 1149 111
rect 1105 74 1107 89
rect 1217 109 1219 112
rect 1147 73 1149 88
rect 1183 83 1185 97
rect 1599 109 1601 112
rect 1217 74 1219 89
rect 1332 76 1334 97
rect 1366 77 1368 97
rect 1413 91 1415 94
rect 654 59 656 63
rect 612 51 614 59
rect 724 51 726 59
rect 851 51 853 60
rect 920 56 922 71
rect 1036 68 1038 72
rect 1530 82 1532 97
rect 1565 83 1567 97
rect 1641 108 1643 111
rect 1599 74 1601 89
rect 1711 109 1713 112
rect 1641 73 1643 88
rect 1677 83 1679 97
rect 1711 74 1713 89
rect 1826 76 1828 97
rect 1860 77 1862 97
rect 1907 91 1909 94
rect 1147 59 1149 63
rect 578 43 580 51
rect 690 43 692 51
rect 612 37 614 41
rect 1105 51 1107 59
rect 1217 51 1219 59
rect 1344 51 1346 60
rect 1413 56 1415 71
rect 1530 68 1532 72
rect 1641 59 1643 63
rect 920 42 922 46
rect 1071 43 1073 51
rect 724 37 726 41
rect 851 37 853 41
rect 1183 43 1185 51
rect 1105 37 1107 41
rect 1599 51 1601 59
rect 1711 51 1713 59
rect 1838 51 1840 60
rect 1907 56 1909 71
rect 1413 42 1415 46
rect 1565 43 1567 51
rect 1217 37 1219 41
rect 1344 37 1346 41
rect 1677 43 1679 51
rect 1599 37 1601 41
rect 1907 42 1909 46
rect 1711 37 1713 41
rect 1838 37 1840 41
rect 578 29 580 33
rect 690 29 692 33
rect 1071 29 1073 33
rect 1183 29 1185 33
rect 1565 29 1567 33
rect 1677 29 1679 33
rect 842 20 844 29
rect 1335 20 1337 29
rect 1829 20 1831 29
rect 842 6 844 10
rect 1335 6 1337 10
rect 1829 6 1831 10
<< polycontact >>
rect 537 85 543 90
rect 572 85 578 90
rect 606 76 612 81
rect 648 76 654 81
rect 684 85 690 90
rect 718 76 724 81
rect 833 78 839 83
rect 875 78 881 83
rect 1030 85 1036 90
rect 1065 85 1071 90
rect 1099 76 1105 81
rect 1141 76 1147 81
rect 1177 85 1183 90
rect 1211 76 1217 81
rect 1326 78 1332 83
rect 1368 78 1374 83
rect 606 54 612 59
rect 718 54 724 59
rect 845 54 851 59
rect 914 59 920 64
rect 1524 85 1530 90
rect 1559 85 1565 90
rect 1593 76 1599 81
rect 1635 76 1641 81
rect 1671 85 1677 90
rect 1705 76 1711 81
rect 1820 78 1826 83
rect 1862 78 1868 83
rect 572 46 578 51
rect 684 46 690 51
rect 1099 54 1105 59
rect 1211 54 1217 59
rect 1338 54 1344 59
rect 1407 59 1413 64
rect 1065 46 1071 51
rect 1177 46 1183 51
rect 1593 54 1599 59
rect 1705 54 1711 59
rect 1832 54 1838 59
rect 1901 59 1907 64
rect 1559 46 1565 51
rect 1671 46 1677 51
rect 836 23 842 28
rect 1329 23 1335 28
rect 1823 23 1829 28
<< metal1 >>
rect 113 171 122 205
rect 0 46 8 162
rect 135 151 144 206
rect 608 172 616 205
rect 12 85 20 142
rect 272 -34 280 69
rect 293 23 301 162
rect 314 61 322 142
rect 465 -34 473 64
rect 494 51 502 162
rect 629 151 637 205
rect 1101 172 1109 205
rect 505 90 513 141
rect 538 122 698 128
rect 537 117 542 122
rect 572 117 577 122
rect 641 119 645 122
rect 546 90 551 97
rect 641 113 669 119
rect 684 117 689 122
rect 586 97 606 104
rect 559 90 564 95
rect 505 85 529 90
rect 534 85 537 90
rect 546 85 572 90
rect 517 59 522 85
rect 546 82 551 85
rect 599 76 606 81
rect 537 67 542 72
rect 615 69 620 89
rect 648 108 653 113
rect 698 97 718 104
rect 657 81 662 88
rect 682 85 684 90
rect 641 76 648 81
rect 657 76 718 81
rect 657 73 662 76
rect 530 62 546 67
rect 551 62 558 67
rect 517 54 606 59
rect 615 51 620 63
rect 648 57 653 63
rect 641 53 669 57
rect 494 46 560 51
rect 566 46 572 51
rect 581 43 606 47
rect 546 5 551 36
rect 572 5 577 33
rect 648 5 653 53
rect 672 51 675 76
rect 727 69 732 89
rect 732 63 774 69
rect 713 54 718 59
rect 727 51 732 63
rect 672 46 684 51
rect 693 43 718 47
rect 684 5 689 33
rect 551 0 700 5
rect 767 -34 774 63
rect 787 28 795 162
rect 808 67 816 141
rect 833 122 904 128
rect 833 117 838 122
rect 867 117 872 122
rect 908 102 913 122
rect 842 83 847 97
rect 876 92 881 97
rect 907 96 935 102
rect 867 88 881 92
rect 914 91 919 96
rect 867 83 872 88
rect 821 78 833 83
rect 842 78 872 83
rect 881 78 886 83
rect 821 67 826 78
rect 808 61 826 67
rect 821 59 826 61
rect 854 64 859 78
rect 923 64 928 71
rect 854 59 914 64
rect 923 59 967 64
rect 821 54 845 59
rect 854 51 859 59
rect 923 56 928 59
rect 787 23 820 28
rect 827 23 836 28
rect 845 20 850 41
rect 914 40 919 46
rect 907 36 935 40
rect 836 4 841 10
rect 912 4 919 36
rect 834 -1 912 4
rect 960 -34 967 59
rect 987 51 995 162
rect 1122 151 1130 205
rect 1595 172 1603 205
rect 998 90 1006 141
rect 1032 122 1191 128
rect 1030 117 1035 122
rect 1065 117 1070 122
rect 1134 119 1138 122
rect 1039 90 1044 97
rect 1134 113 1162 119
rect 1177 117 1182 122
rect 1079 97 1099 104
rect 1052 90 1057 95
rect 998 85 1022 90
rect 1027 85 1030 90
rect 1039 85 1065 90
rect 1010 59 1015 85
rect 1039 82 1044 85
rect 1092 76 1099 81
rect 1030 67 1035 72
rect 1108 69 1113 89
rect 1141 108 1146 113
rect 1191 97 1211 104
rect 1150 81 1155 88
rect 1175 85 1177 90
rect 1134 76 1141 81
rect 1150 76 1211 81
rect 1150 73 1155 76
rect 1023 62 1039 67
rect 1044 62 1051 67
rect 1010 54 1099 59
rect 1108 51 1113 63
rect 1141 57 1146 63
rect 1134 53 1162 57
rect 987 46 1053 51
rect 1059 46 1065 51
rect 1074 43 1099 47
rect 1039 5 1044 36
rect 1065 5 1070 33
rect 1141 5 1146 53
rect 1165 51 1168 76
rect 1220 69 1225 89
rect 1225 63 1267 69
rect 1206 54 1211 59
rect 1220 51 1225 63
rect 1165 46 1177 51
rect 1186 43 1211 47
rect 1177 5 1182 33
rect 1046 0 1192 5
rect 1260 -34 1267 63
rect 1280 28 1288 162
rect 1301 67 1309 141
rect 1326 122 1397 128
rect 1326 117 1331 122
rect 1360 117 1365 122
rect 1401 102 1406 122
rect 1335 83 1340 97
rect 1369 92 1374 97
rect 1400 96 1428 102
rect 1360 88 1374 92
rect 1407 91 1412 96
rect 1360 83 1365 88
rect 1314 78 1326 83
rect 1335 78 1365 83
rect 1374 78 1379 83
rect 1314 67 1319 78
rect 1301 61 1319 67
rect 1314 59 1319 61
rect 1347 64 1352 78
rect 1416 64 1421 71
rect 1347 59 1407 64
rect 1416 59 1460 64
rect 1314 54 1338 59
rect 1347 51 1352 59
rect 1416 56 1421 59
rect 1280 23 1313 28
rect 1320 23 1329 28
rect 1338 20 1343 41
rect 1407 40 1412 46
rect 1400 36 1428 40
rect 1329 4 1334 10
rect 1405 4 1412 36
rect 1328 -1 1407 4
rect 1453 -34 1460 59
rect 1481 51 1489 162
rect 1616 151 1624 205
rect 1492 90 1500 141
rect 1526 122 1685 128
rect 1524 117 1529 122
rect 1559 117 1564 122
rect 1628 119 1632 122
rect 1533 90 1538 97
rect 1628 113 1656 119
rect 1671 117 1676 122
rect 1573 97 1593 104
rect 1546 90 1551 95
rect 1492 85 1516 90
rect 1521 85 1524 90
rect 1533 85 1559 90
rect 1504 59 1509 85
rect 1533 82 1538 85
rect 1586 76 1593 81
rect 1524 67 1529 72
rect 1602 69 1607 89
rect 1635 108 1640 113
rect 1685 97 1705 104
rect 1644 81 1649 88
rect 1669 85 1671 90
rect 1628 76 1635 81
rect 1644 76 1705 81
rect 1644 73 1649 76
rect 1517 62 1533 67
rect 1538 62 1545 67
rect 1504 54 1593 59
rect 1602 51 1607 63
rect 1635 57 1640 63
rect 1628 53 1656 57
rect 1481 46 1547 51
rect 1553 46 1559 51
rect 1568 43 1593 47
rect 1533 5 1538 36
rect 1559 5 1564 33
rect 1635 5 1640 53
rect 1659 51 1662 76
rect 1714 69 1719 89
rect 1719 63 1761 69
rect 1700 54 1705 59
rect 1714 51 1719 63
rect 1659 46 1671 51
rect 1680 43 1705 47
rect 1671 5 1676 33
rect 1538 0 1685 5
rect 1754 -34 1761 63
rect 1774 28 1782 162
rect 1795 67 1803 141
rect 1820 122 1900 128
rect 1820 117 1825 122
rect 1854 117 1859 122
rect 1895 102 1900 122
rect 1829 83 1834 97
rect 1863 92 1868 97
rect 1894 96 1922 102
rect 1854 88 1868 92
rect 1901 91 1906 96
rect 1854 83 1859 88
rect 1808 78 1820 83
rect 1829 78 1859 83
rect 1868 78 1873 83
rect 1808 67 1813 78
rect 1795 61 1813 67
rect 1808 59 1813 61
rect 1841 64 1846 78
rect 1910 64 1915 71
rect 1841 59 1901 64
rect 1910 59 1954 64
rect 1808 54 1832 59
rect 1841 51 1846 59
rect 1910 56 1915 59
rect 1774 23 1807 28
rect 1814 23 1823 28
rect 1832 20 1837 41
rect 1901 40 1906 46
rect 1894 36 1922 40
rect 1823 4 1828 10
rect 1899 4 1906 36
rect 1823 -1 1906 4
rect 1947 -34 1954 59
<< m2contact >>
rect 0 162 8 171
rect 113 162 124 171
rect 293 162 301 171
rect 11 142 20 151
rect 135 142 145 151
rect 204 122 211 128
rect 203 0 211 5
rect 494 162 502 171
rect 608 162 616 172
rect 313 142 322 151
rect 332 122 339 128
rect 412 122 419 128
rect 335 0 343 5
rect 418 0 425 5
rect 505 141 513 150
rect 629 141 637 151
rect 787 162 795 171
rect 529 122 538 128
rect 698 122 705 129
rect 559 95 564 100
rect 529 85 534 90
rect 594 76 599 81
rect 677 85 682 90
rect 636 76 641 81
rect 546 62 551 67
rect 615 63 620 69
rect 560 46 566 51
rect 546 36 551 41
rect 727 63 732 69
rect 706 54 713 59
rect 546 0 551 5
rect 700 0 705 5
rect 987 162 995 171
rect 1101 162 1109 172
rect 808 141 816 150
rect 826 122 833 129
rect 904 122 913 128
rect 886 78 893 83
rect 820 23 827 28
rect 829 -1 834 4
rect 912 -1 919 4
rect 998 141 1006 150
rect 1122 141 1130 151
rect 1280 162 1288 171
rect 1023 122 1032 128
rect 1191 122 1198 129
rect 1052 95 1057 100
rect 1022 85 1027 90
rect 1087 76 1092 81
rect 1170 85 1175 90
rect 1129 76 1134 81
rect 1039 62 1044 67
rect 1108 63 1113 69
rect 1053 46 1059 51
rect 1039 36 1044 41
rect 1220 63 1225 69
rect 1199 54 1206 59
rect 1039 0 1046 5
rect 1192 0 1198 5
rect 1481 162 1489 171
rect 1595 162 1603 172
rect 1301 141 1309 150
rect 1319 122 1326 129
rect 1397 122 1406 128
rect 1379 78 1386 83
rect 1313 23 1320 28
rect 1322 -1 1328 4
rect 1407 -1 1412 4
rect 1492 141 1500 150
rect 1616 141 1624 151
rect 1774 162 1782 171
rect 1517 122 1526 128
rect 1685 122 1692 129
rect 1546 95 1551 100
rect 1516 85 1521 90
rect 1581 76 1586 81
rect 1664 85 1669 90
rect 1623 76 1628 81
rect 1533 62 1538 67
rect 1602 63 1607 69
rect 1547 46 1553 51
rect 1533 36 1538 41
rect 1714 63 1719 69
rect 1693 54 1700 59
rect 1533 0 1538 5
rect 1685 0 1692 5
rect 1795 141 1803 150
rect 1813 122 1820 129
rect 1873 78 1880 83
rect 1807 23 1814 28
rect 1816 -1 1823 4
<< metal2 >>
rect 8 162 113 171
rect 124 162 293 171
rect 502 162 608 171
rect 616 162 787 171
rect 995 162 1101 171
rect 1109 162 1280 171
rect 1489 162 1595 171
rect 1603 162 1774 171
rect 20 142 135 151
rect 145 142 313 151
rect 513 141 629 150
rect 637 141 808 150
rect 1006 141 1122 150
rect 1130 141 1301 150
rect 1500 141 1616 150
rect 1624 141 1795 150
rect 211 122 332 128
rect 419 122 529 128
rect 705 122 826 129
rect 913 122 1023 128
rect 1198 122 1319 129
rect 1406 122 1517 128
rect 1692 122 1813 129
rect 564 95 749 100
rect 1057 95 1242 100
rect 1551 95 1736 100
rect 534 85 677 90
rect 560 76 594 81
rect 599 76 636 81
rect 546 41 551 62
rect 560 51 566 76
rect 620 63 727 69
rect 743 59 749 95
rect 1027 85 1170 90
rect 713 54 749 59
rect 886 28 893 78
rect 1053 76 1087 81
rect 1092 76 1129 81
rect 1039 41 1044 62
rect 1053 51 1059 76
rect 1113 63 1220 69
rect 1236 59 1242 95
rect 1521 85 1664 90
rect 1206 54 1242 59
rect 1379 28 1386 78
rect 1547 76 1581 81
rect 1586 76 1623 81
rect 1533 41 1538 62
rect 1547 51 1553 76
rect 1607 63 1714 69
rect 1730 59 1736 95
rect 1700 54 1736 59
rect 1873 28 1880 78
rect 827 23 893 28
rect 1320 23 1386 28
rect 1814 23 1880 28
rect 211 0 335 5
rect 425 0 546 4
rect 705 0 829 4
rect 418 -1 551 0
rect 919 0 1039 4
rect 1198 0 1322 4
rect 1412 0 1533 4
rect 1692 0 1816 4
rect 1412 -1 1538 0
use xorgate  xorgate_0
timestamp 1618846832
transform 1 0 142 0 1 53
box -142 -53 138 75
use andgate  andgate_0
timestamp 1618846967
transform 1 0 408 0 1 36
box -115 -36 65 92
<< end >>
