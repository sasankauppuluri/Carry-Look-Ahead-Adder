magic
tech scmos
timestamp 1619553084
<< metal1 >>
rect -634 1945 -329 1951
rect 1094 1810 1356 1816
rect 1459 1810 1721 1816
rect -489 1770 -449 1775
rect -80 1770 -39 1776
rect -801 1516 -697 1521
rect -457 1489 -449 1770
rect -46 1629 -39 1770
rect 1241 1635 1271 1640
rect 1605 1635 1635 1640
rect 1964 1635 1994 1640
rect -46 1622 40 1629
rect -8 1596 25 1603
rect -392 1516 -288 1521
rect 0 1489 10 1596
rect -457 1488 -293 1489
rect -142 1488 10 1489
rect -457 1481 10 1488
rect 819 1386 829 1442
rect 819 1381 948 1386
rect 1293 1348 1302 1386
rect 819 1340 1302 1348
rect 819 1323 829 1340
rect 801 1317 829 1323
rect 1652 1320 1663 1386
rect 878 1310 1663 1320
rect -489 1279 -449 1284
rect -80 1279 -39 1284
rect -801 1025 -697 1030
rect -457 994 -449 1279
rect -46 1137 -39 1279
rect 878 1181 890 1310
rect 816 1175 890 1181
rect -46 1130 40 1137
rect 1241 1124 1271 1129
rect 1605 1124 1635 1129
rect 0 1112 9 1113
rect -8 1105 25 1112
rect -392 1025 -288 1030
rect 0 994 9 1105
rect 858 1039 865 1040
rect 826 1033 865 1039
rect -457 986 9 994
rect -457 985 -449 986
rect 818 891 837 897
rect 830 840 837 891
rect 858 875 865 1033
rect 858 870 937 875
rect 1293 840 1299 875
rect 830 833 1299 840
rect -489 789 -449 794
rect -59 789 -39 794
rect -801 535 -697 540
rect -457 506 -449 789
rect -69 666 -62 671
rect -45 646 -39 789
rect -45 639 40 646
rect -8 614 25 621
rect -392 535 -288 540
rect 0 506 9 614
rect 1899 580 1929 585
rect -457 498 9 506
rect 1911 392 1941 397
rect -461 298 -449 303
rect -51 298 -39 303
rect -802 44 -697 49
rect -457 13 -449 298
rect -45 155 -39 298
rect 1929 204 1959 209
rect -45 148 40 155
rect -9 123 25 130
rect -392 44 -288 49
rect -1 13 10 123
rect 1946 42 1977 49
rect 360 24 374 30
rect -457 5 10 13
<< m2contact >>
rect -784 1647 -778 1652
rect -375 1647 -369 1652
rect 945 1512 954 1517
rect 1307 1512 1314 1517
rect 1666 1512 1673 1517
rect -784 1156 -778 1161
rect -374 1156 -368 1161
rect 946 1001 954 1006
rect 1307 1001 1314 1006
rect 1162 845 1170 851
rect 1401 846 1409 851
rect -784 666 -778 671
rect -374 666 -368 671
rect -784 175 -778 180
rect -568 19 -560 25
rect -375 175 -369 180
rect -284 20 -277 25
<< metal2 >>
rect -583 1964 -565 2003
rect -784 1957 953 1964
rect -784 1652 -778 1957
rect -784 1161 -778 1647
rect -375 1652 -369 1957
rect -745 1454 -738 1592
rect -784 671 -778 1156
rect -375 1161 -369 1647
rect 946 1832 953 1957
rect 946 1823 1673 1832
rect -336 1454 -329 1592
rect 946 1517 953 1823
rect 1307 1517 1314 1823
rect -375 1156 -374 1161
rect -745 964 -738 1102
rect -784 180 -778 666
rect -375 671 -369 1156
rect -336 964 -329 1102
rect 946 1006 954 1512
rect 1666 1517 1673 1823
rect 985 1299 992 1457
rect 1307 1006 1314 1512
rect 1349 1299 1356 1457
rect 946 1000 954 1001
rect 1170 846 1401 851
rect 1170 845 1409 846
rect -375 666 -374 671
rect -745 473 -738 611
rect -375 180 -369 666
rect -336 473 -329 611
rect -560 20 -284 25
rect -560 19 -277 20
<< m123contact >>
rect 1760 1357 1767 1362
<< metal3 >>
rect -504 1360 -497 1623
rect -95 1360 -88 1623
rect 1226 1205 1233 1488
rect 1590 1362 1597 1488
rect 1590 1357 1760 1362
rect 1590 1205 1597 1357
rect -504 870 -497 1133
rect -95 869 -88 1132
rect -504 379 -497 642
rect -95 379 -88 642
use dff  dff_7
timestamp 1619529728
transform 1 0 -587 0 1 1741
box -214 -250 128 210
use dff  dff_6
timestamp 1619529728
transform 1 0 -178 0 1 1741
box -214 -250 128 210
use dff  dff_5
timestamp 1619529728
transform 1 0 -587 0 1 1250
box -214 -250 128 210
use dff  dff_4
timestamp 1619529728
transform 1 0 -178 0 1 1250
box -214 -250 128 210
use dff  dff_10
timestamp 1619529728
transform 1 0 1143 0 1 1606
box -214 -250 128 210
use dff  dff_11
timestamp 1619529728
transform 1 0 1507 0 1 1606
box -214 -250 128 210
use dff  dff_12
timestamp 1619529728
transform 1 0 1866 0 1 1606
box -214 -250 128 210
use dff  dff_3
timestamp 1619529728
transform 1 0 -587 0 1 760
box -214 -250 128 210
use dff  dff_2
timestamp 1619529728
transform 1 0 -178 0 1 760
box -214 -250 128 210
use dff  dff_8
timestamp 1619529728
transform 1 0 1143 0 1 1095
box -214 -250 128 210
use dff  dff_9
timestamp 1619529728
transform 1 0 1507 0 1 1095
box -214 -250 128 210
use dff  dff_1
timestamp 1619529728
transform 1 0 -587 0 1 269
box -214 -250 128 210
use dff  dff_0
timestamp 1619529728
transform 1 0 -178 0 1 269
box -214 -250 128 210
use clablock  clablock_0
timestamp 1619544759
transform 1 0 -8 0 1 5
box 0 -5 1998 1942
<< labels >>
rlabel metal2 -583 1964 -566 2003 1 clk
rlabel space 176 -213 279 -109 1 DA0
rlabel metal1 -802 44 -697 49 1 DA0
rlabel metal1 -801 535 -697 540 1 DA1
rlabel metal1 -801 1025 -697 1030 1 DA2
rlabel metal1 -801 1516 -697 1521 1 DA3
rlabel metal1 -392 1516 -288 1521 1 DB3
rlabel metal1 -392 1025 -288 1030 1 DB2
rlabel metal1 -392 535 -288 540 1 DB1
rlabel metal1 -392 44 -288 49 1 DB0
rlabel metal1 -9 123 25 130 1 A0
rlabel metal1 -8 614 25 621 1 A1
rlabel metal1 -8 1105 25 1112 1 A2
rlabel metal1 -8 1596 25 1603 1 A3
rlabel metal1 -8 1622 40 1629 1 B3
rlabel metal1 -8 1130 40 1137 1 B2
rlabel metal1 -8 639 40 646 1 B1
rlabel metal1 -9 148 40 155 1 B0
rlabel metal1 360 24 374 30 1 Car0
rlabel metal1 1946 42 1977 49 1 Car1
rlabel metal1 1929 204 1959 209 1 Car2
rlabel metal1 1911 392 1941 397 1 Car3
rlabel metal1 818 891 837 897 1 S0
rlabel metal1 837 1033 865 1039 1 S1
rlabel metal1 837 1175 865 1181 1 S2
rlabel metal1 801 1317 829 1323 1 S3
rlabel metal1 1899 580 1929 585 1 Carout
rlabel metal1 1605 1124 1635 1129 1 Q0
rlabel metal1 1241 1124 1271 1129 1 Q1
rlabel metal1 1964 1635 1994 1640 1 Q2
rlabel metal1 1605 1635 1635 1640 1 Q3
rlabel metal1 1241 1635 1271 1640 1 Q4
<< end >>
